// Copyright (c) UnnamedOrange and Jack-Lyu. Licensed under the MIT License.
// See the LICENSE file in the repository root for full license text.

/// <projectname>mania-to-go</projectname>
/// <modulename>update_others_t</modulename>
/// <filedescription>update ������Ϣ������ʱ�䡢���ء��ܷ�����</filedescription>
/// <version>
/// 0.0.1 (UnnamedOrange) : First commit.
/// </version>

`timescale 1ns / 1ps

module update_others_t #
(
	// �ڲ�������
	parameter state_width = 4
)
(
	// ���ơ�
	input sig_on,
	output sig_done,

	// BRAM��
	output reg [11:0] dt_b_addr,
	input [31:0] dt_b_data_out,
	output reg dt_b_en,

	// ���������ַ��
	input [11:0] dt_size,
	input [11:0] dt_base_addr, // == 2

	// ��Ϸ״̬��
	input [3:0] is_game_over,
	input [7:0] is_combo,
	input [3:0] is_miss,
	input [3:0] is_bad,
	input [3:0] is_good,
	input [3:0] is_great,
	input [3:0] is_perfect,
	input [19:0] song_length,

	// ��Ҫ��Ϊ����ı�����
	output reg [19:0] current_time,
	output reg [31:0] current_pixel,

	output reg [15:0] miss,
	output reg [15:0] bad,
	output reg [15:0] good,
	output reg [15:0] great,
	output reg [15:0] perfect,
	output reg [15:0] combo,

	output reg [3:0] current_score, // 0 Ϊ�գ�Ȼ�������� perfect, great, good, bad, miss��
	output reg [1:0] current_score_fade,

	// ��λ��ʱ�ӡ�
	input RESET_L,
	input CLK
);

	// ������
	reg [11:0] current_speed;
	reg [11:0] current_offset;

	// ״̬���塣
	localparam [state_width - 1 : 0]
		s_init                     = 4'd0,       // ��λ��
		s_update_speed             = 4'd1,       // �����ٶȡ�
		s_w_update_speed           = 4'd2,       // �ȴ������ٶȡ�
		s_update_time_and_pixel    = 4'd3,       // ����ʱ������ء�
		s_update_score             = 4'd4,       // ���·�����
		s_done                     = 4'b1111,    // ��ɡ�
		s_unused = 4'b1111;
	reg [state_width - 1 : 0] state, n_state;

	// ��ȡ�������ٶȡ�
	wire sig_update_speed_on;
	reg sig_update_speed_done;
	always @(posedge CLK) begin : update_speed_t
		reg working;
		reg [1:0] pat;

		if (!RESET_L) begin
			current_speed <= 0;
			current_offset <= 0;
			working <= 0;
			pat <= 0;
			sig_update_speed_done <= 0;
			dt_b_addr <= 0;
			dt_b_en <= 0;
		end
		else begin
			if (!working) begin
				if (sig_update_speed_on)
					working <= 1;
			end
			else begin
				if (pat == 0) begin
					dt_b_en <= 1;
					dt_b_addr <= dt_base_addr + current_offset;
				end
				else if (pat == 3) begin
					dt_b_en <= 0;
					working <= 0;
					// �����ٶȡ�
					if (dt_b_data_out[19:0] == current_time) begin
						current_speed <= dt_b_data_out[31:20];
						current_offset <= current_offset + 1;
					end
				end
				pat <= pat + 1;
			end
			sig_update_speed_done <= working && pat == 2'b11;
		end
	end

	// ����ʱ���λ�á�
	always @(posedge CLK) begin
		if (!RESET_L) begin
			current_time <= 0;
			current_pixel <= 0;
		end
		else begin
			if (state == s_update_time_and_pixel) begin
				if (current_time < song_length) begin
					current_time <= current_time + 1;
					current_pixel <= current_pixel + current_speed;
				end
			end
		end
	end

	// ���·�����
	reg [15:0] next_miss;
	reg [15:0] next_bad;
	reg [15:0] next_good;
	reg [15:0] next_great;
	reg [15:0] next_perfect;
	reg [15:0] next_combo;
	reg [3:0] next_current_score;
	reg [15:0] score_counter;
	reg [15:0] next_score_counter;
	parameter fade_time = 350;
	always @(posedge CLK) begin
		if (!RESET_L) begin
			miss <= 0;
			bad <= 0;
			good <= 0;
			great <= 0;
			perfect <= 0;
			combo <= 0;
			current_score <= 0;
			score_counter <= 0;
		end
		else begin
			if (state == s_update_score) begin
				miss <= next_miss;
				bad <= next_bad;
				good <= next_good;
				great <= next_great;
				perfect <= next_perfect;
				combo <= next_combo;
				current_score <= next_current_score;
				score_counter <= next_score_counter;
			end
		end
	end

	always @(*) begin : score_excitation
		integer i, j;

		next_miss = miss;
		next_bad = bad;
		next_good = good;
		next_great = great;
		next_perfect = perfect;
		for (i = 0; i < 4; i = i + 1) begin
			next_miss = next_miss + is_miss[i];
			for (j = 0; j < 4; j = j + 1) begin
				if (next_miss[j * 4 +: 4] >= 10) begin
					next_miss[j * 4 +: 4] = 0;
					if (j + 1 < 4)
						next_miss[(j + 1) * 4 +: 4] = next_miss[(j + 1) * 4 +: 4] + 1;
				end
			end
		end
		for (i = 0; i < 4; i = i + 1) begin
			next_bad = next_bad + is_bad[i];
			for (j = 0; j < 4; j = j + 1) begin
				if (next_bad[j * 4 +: 4] >= 10) begin
					next_bad[j * 4 +: 4] = 0;
					if (j + 1 < 4)
						next_bad[(j + 1) * 4 +: 4] = next_bad[(j + 1) * 4 +: 4] + 1;
				end
			end
		end
		for (i = 0; i < 4; i = i + 1) begin
			next_good = next_good + is_good[i];
			for (j = 0; j < 4; j = j + 1) begin
				if (next_good[j * 4 +: 4] >= 10) begin
					next_good[j * 4 +: 4] = 0;
					if (j + 1 < 4)
						next_good[(j + 1) * 4 +: 4] = next_good[(j + 1) * 4 +: 4] + 1;
				end
			end
		end
		for (i = 0; i < 4; i = i + 1) begin
			next_great = next_great + is_great[i];
			for (j = 0; j < 4; j = j + 1) begin
				if (next_great[j * 4 +: 4] >= 10) begin
					next_great[j * 4 +: 4] = 0;
					if (j + 1 < 4)
						next_great[(j + 1) * 4 +: 4] = next_great[(j + 1) * 4 +: 4] + 1;
				end
			end
		end
		for (i = 0; i < 4; i = i + 1) begin
			next_perfect = next_perfect + is_perfect[i];
			for (j = 0; j < 4; j = j + 1) begin
				if (next_perfect[j * 4 +: 4] >= 10) begin
					next_perfect[j * 4 +: 4] = 0;
					if (j + 1 < 4)
						next_perfect[(j + 1) * 4 +: 4] = next_perfect[(j + 1) * 4 +: 4] + 1;
				end
			end
		end

		next_combo = combo;
		for (i = 0; i < 4; i = i + 1)
			if (is_combo[i * 2 +: 2] == 2'b10)
				next_combo = 0;
		for (i = 0; i < 4; i = i + 1) begin
			if (is_combo[i * 2 +: 2] == 2'b01)
				next_combo = next_combo + 1;
			for (j = 0; j < 4; j = j + 1) begin
				if (next_combo[j * 4 +: 4] >= 10) begin
					next_combo[j * 4 +: 4] = 0;
					if (j + 1 < 4)
						next_combo[(j + 1) * 4 +: 4] = next_combo[(j + 1) * 4 +: 4] + 1;
				end
			end
		end

		next_current_score = current_score;
		next_score_counter = score_counter ? score_counter - 1 : 0;
		for (i = 0; i < 4; i = i + 1)
			if (is_perfect[i]) begin
				next_current_score = 1;
				next_score_counter = fade_time;
			end
		for (i = 0; i < 4; i = i + 1)
			if (is_great[i]) begin
				next_current_score = 2;
				next_score_counter = fade_time;
			end
		for (i = 0; i < 4; i = i + 1)
			if (is_good[i]) begin
				next_current_score = 3;
				next_score_counter = fade_time;
			end
		for (i = 0; i < 4; i = i + 1)
			if (is_bad[i]) begin
				next_current_score = 4;
				next_score_counter = fade_time;
			end
		for (i = 0; i < 4; i = i + 1)
			if (is_miss[i]) begin
				next_current_score = 5;
				next_score_counter = fade_time;
			end
		if (next_score_counter == 0)
			next_current_score = 0;
	end

	always @(*) begin
		if (score_counter == 0)
			current_score_fade = 0;
		if (score_counter < 30)
			current_score_fade = 3;
		else if (score_counter < 60)
			current_score_fade = 2;
		else if (score_counter < fade_time - 30)
			current_score_fade = 0;
		else
			current_score_fade = 1;
	end

	// �������̡�
	always @(posedge CLK) begin
		if (!RESET_L) begin
			state <= s_init;
		end
		else begin
			state <= n_state;
		end
	end

	// �������̡�
	always @(*) begin
		case (state)
			s_init:
				n_state = sig_on ? ((current_offset < dt_size) ? s_update_speed : s_update_time_and_pixel) : s_init;
			s_update_speed:
				n_state = s_w_update_speed;
			s_w_update_speed:
				n_state = sig_update_speed_done ? s_update_time_and_pixel : s_w_update_speed;
			s_update_time_and_pixel:
				n_state = s_update_score;
			s_update_score:
				n_state = s_done;
			s_done:
				n_state = s_init;
			default:
				n_state = s_init;
		endcase
	end

	// ������̡�
	assign sig_done = state == s_done;
	assign sig_update_speed_on = state == s_update_speed;

endmodule